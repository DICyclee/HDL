/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2024 Spring ---------------------- //
// ---------------------- Editor : 	David   -----------------------//
// ---------------------- Date : 2024.01    ---------------------- //
// ----------------------      test1        ---------------------- //
// --------------------  Bitwise operator  ------------------------//
/////////////////////////////////////////////////////////////////////
module test1(out1, 
             out2,
             out3,
             out4,
             in1, 
             in2);
             
input  [2:0] in1,  in2;
output [2:0] out1, out2, out3, out4;
	
assign out1 = in1 & in2;  //and
assign out2 = in1 | in2;  //or
assign out3 = in1 ^ in2;  //xor
assign out4 = ~in1;       //not
	
endmodule